module initial_bad();
reg clk,reset;
wire enable,data;

initial begin
 clk = 0;
 reset = 0;
 enable = 0;
 data = 0;
end

endmodule
